module BUF(in,out);
input in;
output out;
assign #5 out=in;
endmodule